-- SIPO (Serial-In Parallel-Out) Register
-- By: Ryan Vickramasinghe